
module color_map
(
    input [7:0] value,
    output reg [23:0] rgb
);
    always @(*) begin
        case (value)

             8'd0   : rgb = 24'hff6666;
             8'd128 : rgb = 24'hcd3434;
             8'd1   : rgb = 24'hff6d66;
             8'd129 : rgb = 24'hcd3b34;
             8'd2   : rgb = 24'hff7466;
             8'd130 : rgb = 24'hcd4234;
             8'd3   : rgb = 24'hff7c66;
             8'd131 : rgb = 24'hcd4a34;
             8'd4   : rgb = 24'hff8366;
             8'd132 : rgb = 24'hcd5134;
             8'd5   : rgb = 24'hff8a66;
             8'd133 : rgb = 24'hcd5834;
             8'd6   : rgb = 24'hff9166;
             8'd134 : rgb = 24'hcd5f34;
             8'd7   : rgb = 24'hff9866;
             8'd135 : rgb = 24'hcd6634;
             8'd8   : rgb = 24'hff9f66;
             8'd136 : rgb = 24'hcd6d34;
             8'd9   : rgb = 24'hffa766;
             8'd137 : rgb = 24'hcd7534;
             8'd10  : rgb = 24'hffae66;
             8'd138 : rgb = 24'hcd7c34;
             8'd11  : rgb = 24'hffb566;
             8'd139 : rgb = 24'hcd8334;
             8'd12  : rgb = 24'hffbc66;
             8'd140 : rgb = 24'hcd8a34;
             8'd13  : rgb = 24'hffc366;
             8'd141 : rgb = 24'hcd9134;
             8'd14  : rgb = 24'hffca66;
             8'd142 : rgb = 24'hcd9834;
             8'd15  : rgb = 24'hffd266;
             8'd143 : rgb = 24'hcda034;
             8'd16  : rgb = 24'hffd966;
             8'd144 : rgb = 24'hcda734;
             8'd17  : rgb = 24'hffe066;
             8'd145 : rgb = 24'hcdae34;
             8'd18  : rgb = 24'hffe766;
             8'd146 : rgb = 24'hcdb534;
             8'd19  : rgb = 24'hffee66;
             8'd147 : rgb = 24'hcdbc34;
             8'd20  : rgb = 24'hfff566;
             8'd148 : rgb = 24'hcdc334;
             8'd21  : rgb = 24'hfffd66;
             8'd149 : rgb = 24'hcdcb34;
             8'd22  : rgb = 24'hfaff66;
             8'd150 : rgb = 24'hc8cd34;
             8'd23  : rgb = 24'hf3ff66;
             8'd151 : rgb = 24'hc1cd34;
             8'd24  : rgb = 24'hecff66;
             8'd152 : rgb = 24'hbacd34;
             8'd25  : rgb = 24'he5ff66;
             8'd153 : rgb = 24'hb3cd34;
             8'd26  : rgb = 24'hdeff66;
             8'd154 : rgb = 24'haccd34;
             8'd27  : rgb = 24'hd6ff66;
             8'd155 : rgb = 24'ha4cd34;
             8'd28  : rgb = 24'hcfff66;
             8'd156 : rgb = 24'h9dcd34;
             8'd29  : rgb = 24'hc8ff66;
             8'd157 : rgb = 24'h96cd34;
             8'd30  : rgb = 24'hc1ff66;
             8'd158 : rgb = 24'h8fcd34;
             8'd31  : rgb = 24'hbaff66;
             8'd159 : rgb = 24'h88cd34;
             8'd32  : rgb = 24'hb2ff66;
             8'd160 : rgb = 24'h80cd34;
             8'd33  : rgb = 24'habff66;
             8'd161 : rgb = 24'h79cd34;
             8'd34  : rgb = 24'ha4ff66;
             8'd162 : rgb = 24'h72cd34;
             8'd35  : rgb = 24'h9dff66;
             8'd163 : rgb = 24'h6bcd34;
             8'd36  : rgb = 24'h96ff66;
             8'd164 : rgb = 24'h64cd34;
             8'd37  : rgb = 24'h8fff66;
             8'd165 : rgb = 24'h5dcd34;
             8'd38  : rgb = 24'h87ff66;
             8'd166 : rgb = 24'h55cd34;
             8'd39  : rgb = 24'h80ff66;
             8'd167 : rgb = 24'h4ecd34;
             8'd40  : rgb = 24'h79ff66;
             8'd168 : rgb = 24'h47cd34;
             8'd41  : rgb = 24'h72ff66;
             8'd169 : rgb = 24'h40cd34;
             8'd42  : rgb = 24'h6bff66;
             8'd170 : rgb = 24'h39cd34;
             8'd43  : rgb = 24'h66ff68;
             8'd171 : rgb = 24'h34cd36;
             8'd44  : rgb = 24'h66ff70;
             8'd172 : rgb = 24'h34cd3e;
             8'd45  : rgb = 24'h66ff77;
             8'd173 : rgb = 24'h34cd45;
             8'd46  : rgb = 24'h66ff7e;
             8'd174 : rgb = 24'h34cd4c;
             8'd47  : rgb = 24'h66ff85;
             8'd175 : rgb = 24'h34cd53;
             8'd48  : rgb = 24'h66ff8c;
             8'd176 : rgb = 24'h34cd5a;
             8'd49  : rgb = 24'h66ff93;
             8'd177 : rgb = 24'h34cd61;
             8'd50  : rgb = 24'h66ff9b;
             8'd178 : rgb = 24'h34cd69;
             8'd51  : rgb = 24'h66ffa2;
             8'd179 : rgb = 24'h34cd70;
             8'd52  : rgb = 24'h66ffa9;
             8'd180 : rgb = 24'h34cd77;
             8'd53  : rgb = 24'h66ffb0;
             8'd181 : rgb = 24'h34cd7e;
             8'd54  : rgb = 24'h66ffb7;
             8'd182 : rgb = 24'h34cd85;
             8'd55  : rgb = 24'h66ffbe;
             8'd183 : rgb = 24'h34cd8c;
             8'd56  : rgb = 24'h66ffc6;
             8'd184 : rgb = 24'h34cd94;
             8'd57  : rgb = 24'h66ffcd;
             8'd185 : rgb = 24'h34cd9b;
             8'd58  : rgb = 24'h66ffd4;
             8'd186 : rgb = 24'h34cda2;
             8'd59  : rgb = 24'h66ffdb;
             8'd187 : rgb = 24'h34cda9;
             8'd60  : rgb = 24'h66ffe2;
             8'd188 : rgb = 24'h34cdb0;
             8'd61  : rgb = 24'h66ffe9;
             8'd189 : rgb = 24'h34cdb7;
             8'd62  : rgb = 24'h66fff1;
             8'd190 : rgb = 24'h34cdbf;
             8'd63  : rgb = 24'h66fff8;
             8'd191 : rgb = 24'h34cdc6;
             8'd64  : rgb = 24'h66ffff;
             8'd192 : rgb = 24'h34cdcd;
             8'd65  : rgb = 24'h66f8ff;
             8'd193 : rgb = 24'h34c6cd;
             8'd66  : rgb = 24'h66f1ff;
             8'd194 : rgb = 24'h34bfcd;
             8'd67  : rgb = 24'h66e9ff;
             8'd195 : rgb = 24'h34b7cd;
             8'd68  : rgb = 24'h66e2ff;
             8'd196 : rgb = 24'h34b0cd;
             8'd69  : rgb = 24'h66dbff;
             8'd197 : rgb = 24'h34a9cd;
             8'd70  : rgb = 24'h66d4ff;
             8'd198 : rgb = 24'h34a2cd;
             8'd71  : rgb = 24'h66cdff;
             8'd199 : rgb = 24'h349bcd;
             8'd72  : rgb = 24'h66c6ff;
             8'd200 : rgb = 24'h3494cd;
             8'd73  : rgb = 24'h66beff;
             8'd201 : rgb = 24'h348ccd;
             8'd74  : rgb = 24'h66b7ff;
             8'd202 : rgb = 24'h3485cd;
             8'd75  : rgb = 24'h66b0ff;
             8'd203 : rgb = 24'h347ecd;
             8'd76  : rgb = 24'h66a9ff;
             8'd204 : rgb = 24'h3477cd;
             8'd77  : rgb = 24'h66a2ff;
             8'd205 : rgb = 24'h3470cd;
             8'd78  : rgb = 24'h669bff;
             8'd206 : rgb = 24'h3469cd;
             8'd79  : rgb = 24'h6693ff;
             8'd207 : rgb = 24'h3461cd;
             8'd80  : rgb = 24'h668cff;
             8'd208 : rgb = 24'h345acd;
             8'd81  : rgb = 24'h6685ff;
             8'd209 : rgb = 24'h3453cd;
             8'd82  : rgb = 24'h667eff;
             8'd210 : rgb = 24'h344ccd;
             8'd83  : rgb = 24'h6677ff;
             8'd211 : rgb = 24'h3445cd;
             8'd84  : rgb = 24'h6670ff;
             8'd212 : rgb = 24'h343ecd;
             8'd85  : rgb = 24'h6668ff;
             8'd213 : rgb = 24'h3436cd;
             8'd86  : rgb = 24'h6b66ff;
             8'd214 : rgb = 24'h3934cd;
             8'd87  : rgb = 24'h7266ff;
             8'd215 : rgb = 24'h4034cd;
             8'd88  : rgb = 24'h7966ff;
             8'd216 : rgb = 24'h4734cd;
             8'd89  : rgb = 24'h8066ff;
             8'd217 : rgb = 24'h4e34cd;
             8'd90  : rgb = 24'h8766ff;
             8'd218 : rgb = 24'h5534cd;
             8'd91  : rgb = 24'h8f66ff;
             8'd219 : rgb = 24'h5d34cd;
             8'd92  : rgb = 24'h9666ff;
             8'd220 : rgb = 24'h6434cd;
             8'd93  : rgb = 24'h9d66ff;
             8'd221 : rgb = 24'h6b34cd;
             8'd94  : rgb = 24'ha466ff;
             8'd222 : rgb = 24'h7234cd;
             8'd95  : rgb = 24'hab66ff;
             8'd223 : rgb = 24'h7934cd;
             8'd96  : rgb = 24'hb266ff;
             8'd224 : rgb = 24'h8034cd;
             8'd97  : rgb = 24'hba66ff;
             8'd225 : rgb = 24'h8834cd;
             8'd98  : rgb = 24'hc166ff;
             8'd226 : rgb = 24'h8f34cd;
             8'd99  : rgb = 24'hc866ff;
             8'd227 : rgb = 24'h9634cd;
             8'd100 : rgb = 24'hcf66ff;
             8'd228 : rgb = 24'h9d34cd;
             8'd101 : rgb = 24'hd666ff;
             8'd229 : rgb = 24'ha434cd;
             8'd102 : rgb = 24'hde66ff;
             8'd230 : rgb = 24'hac34cd;
             8'd103 : rgb = 24'he566ff;
             8'd231 : rgb = 24'hb334cd;
             8'd104 : rgb = 24'hec66ff;
             8'd232 : rgb = 24'hba34cd;
             8'd105 : rgb = 24'hf366ff;
             8'd233 : rgb = 24'hc134cd;
             8'd106 : rgb = 24'hfa66ff;
             8'd234 : rgb = 24'hc834cd;
             8'd107 : rgb = 24'hff66fd;
             8'd235 : rgb = 24'hcd34cb;
             8'd108 : rgb = 24'hff66f5;
             8'd236 : rgb = 24'hcd34c3;
             8'd109 : rgb = 24'hff66ee;
             8'd237 : rgb = 24'hcd34bc;
             8'd110 : rgb = 24'hff66e7;
             8'd238 : rgb = 24'hcd34b5;
             8'd111 : rgb = 24'hff66e0;
             8'd239 : rgb = 24'hcd34ae;
             8'd112 : rgb = 24'hff66d9;
             8'd240 : rgb = 24'hcd34a7;
             8'd113 : rgb = 24'hff66d2;
             8'd241 : rgb = 24'hcd34a0;
             8'd114 : rgb = 24'hff66ca;
             8'd242 : rgb = 24'hcd3498;
             8'd115 : rgb = 24'hff66c3;
             8'd243 : rgb = 24'hcd3491;
             8'd116 : rgb = 24'hff66bc;
             8'd244 : rgb = 24'hcd348a;
             8'd117 : rgb = 24'hff66b5;
             8'd245 : rgb = 24'hcd3483;
             8'd118 : rgb = 24'hff66ae;
             8'd246 : rgb = 24'hcd347c;
             8'd119 : rgb = 24'hff66a7;
             8'd247 : rgb = 24'hcd3475;
             8'd120 : rgb = 24'hff669f;
             8'd248 : rgb = 24'hcd346d;
             8'd121 : rgb = 24'hff6698;
             8'd249 : rgb = 24'hcd3466;
             8'd122 : rgb = 24'hff6691;
             8'd250 : rgb = 24'hcd345f;
             8'd123 : rgb = 24'hff668a;
             8'd251 : rgb = 24'hcd3458;
             8'd124 : rgb = 24'hff6683;
             8'd252 : rgb = 24'hcd3451;
             8'd125 : rgb = 24'hff667c;
             8'd253 : rgb = 24'hcd344a;
             8'd126 : rgb = 24'hff6674;
             8'd254 : rgb = 24'hcd3442;
             8'd127 : rgb = 24'hff666d;
             8'd255 : rgb = 24'hcd343b;

        endcase
    end
endmodule

