parameter DRAW_MANDELBROT = 2'd0; // Draw binary mandelbrot
parameter DRAW_JULIA = 2'd1;      // Draw julia overlay
parameter DRAW_CLEAR = 2'd2;      // Clear julia overlay
