parameter WRITE_BURST = 1;
parameter READ_BURST_LENGTH = 8;

parameter CMD_IDLE  = 2'd0;
parameter CMD_WRITE = 2'd1;
parameter CMD_READ  = 2'd2;
